*Custom Designer (TM) Version J-2014.12-SP2-2
*Fri Feb  2 04:01:44 2018

*.SCALE METER
*.LDD

********************************************************************************
* Library          : vlsi_lib
* Cell             : nand
* View             : schematic
* View Search List : auCdl schematic symbol
* View Stop List   : auCdl
********************************************************************************
.subckt nand A B VDD VOUT VSS
*.PININFO A:I B:I VDD:I VOUT:O VSS:I
MM5 net21 B VSS VSS n12 w=0.5u l=0.1u nf=1.0 m=1
MM2 VOUT A net21 net21 n12 w=0.5u l=0.1u nf=1.0 m=1
MM4 VOUT A VDD VDD p12 w=0.5u l=0.1u nf=1.0 m=1
MM3 VOUT B VDD net14 p12 w=0.5u l=0.1u nf=1.0 m=1
.ends nand


